package package_comp;
	`include "uvm_macros.svh"
	import  uvm_pkg::*;
	`include "configuration_comp.sv"
	`include "sequencer_comp.sv"	
	`include "driver_comp.sv"
	`include "monitor_comp.sv"
	`include "model_comp.sv"
	`include "agent_comp.sv"
	`include "environment_comp.sv"
	`include "testcase_comp.sv"
endpackage